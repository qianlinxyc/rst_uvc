package rst_uvc_pkg;
    import uvm_pkg::*;

    `include "rst_uvc_cfg.sv"
    `include "rst_uvc_drv.sv"
    `include "rst_uvc_agt.sv"
endpackage : rst_uvc_pkg
